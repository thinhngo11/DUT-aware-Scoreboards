interface my_ifI;
  bit clk, q, qreg;
endinterface
